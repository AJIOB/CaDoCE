library IEEE;
use IEEE.std_logic_1164.all;

entity schema is
  port (
    x1, x2, x3, x4: in std_logic;
    y1, y2, y3, y4: out std_logic
  ) ;
end schema ;

architecture main_arch of schema is

begin

end main_arch ; -- main_arch
